module decodificador (I, O);

	input [3:0] I;
	output reg[6:0] O;

	always @(I) begin
		case (I[3:0])
			'b0000: O = 'b0000001;
			'b0001: O = 'b1001111;
			'b0010: O = 'b0010010;
			'b0011: O = 'b0000110;
			'b0100: O = 'b1001100;
			'b0101: O = 'b0100100;
			'b0110: O = 'b0100000;
			'b0111: O = 'b0001111;
			'b1000: O = 'b0000000;
			'b1001: O = 'b0000100;
			'b1010: O = 'b0001000;
			'b1011: O = 'b1100000;
			'b1100: O = 'b0110001;
			'b1101: O = 'b1000010;
			'b1110: O = 'b0110000;
			'b1111: O = 'b0111000;
		endcase
	end

endmodule 